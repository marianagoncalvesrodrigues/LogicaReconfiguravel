-- Copyright (C) 2019  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
-- Created on Thu Sep 22 11:44:13 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY projeto IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        w : IN STD_LOGIC := '0';
        z : OUT STD_LOGIC;
		  saidaled : OUT STD_LOGIC
    );
END projeto;

ARCHITECTURE BEHAVIOR OF projeto IS
    TYPE type_fstate IS (A,B);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
	 signal ticks: integer:=0;
	 signal cont : integer:=0;
	 constant clockfre: integer := 50e6;
	 
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='0') THEN
            fstate <= A;
        ELSIF rising_edge(clock) THEN
			if ticks = clockfre -1 then
				ticks <= 0;
				saidaled <= '1';
				if cont > 3 then
					cont <= 0;
					saidaled <= '0';
					fstate <= reg_fstate;
				else
					cont <= cont + 1;
				end if;
			else
				ticks <= ticks + 1;
			end if;
				
        END IF;
    END PROCESS;

    PROCESS (fstate,w)
    BEGIN
        z <= '0';
        CASE fstate IS
            WHEN A =>
                IF ((w = '1')) THEN
                    reg_fstate <= B;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= A;
                END IF;
            WHEN B =>
                IF (NOT((w = '1'))) THEN
                    reg_fstate <= A;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= B;
                END IF;

                IF ((w = '1')) THEN
                    z <= '1';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    z <= '0';
                END IF;
            WHEN OTHERS => 
                z <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
